year|indiv|zit|xit
1977|A|1.2|0.6
1977|B|1.5|0.5
1977|C|1.7|0.8
1978|A|0.2|0.06
1978|B|0.7|0.2
1978|C|0.8|0.3
1978|D|0.9|0.5
